//////////////////////////////////////////////////////////////////////////////////////////
//
//  File Name   : ace_dispatch.v
//  Author      : ejune@aureage.com
//                
//  Description : dispatch module dispatches renamed packets to Issue Queue, Active
//                List, and Load-Store queue.
//                Before dipatching it checks if there is enough space for incoming
//                instructions in Issue Queue, Active List, and Load-Store queue.
//                Dispatch width is same as rename width 
//                
//                
//  Create Date : original_time
//  Version     : v0.1 
//
//////////////////////////////////////////////////////////////////////////////////////////
module ace_dispatch ();


endmodule
