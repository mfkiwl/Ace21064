//////////////////////////////////////////////////////////////////////////////////////////
//
//  File Name   : rob.v
//  Author      : ejune@aureage.com
//                
//  Description : reorder buffer is a circular buffer with head and tail pointers. 
//                New instructions are written at tail and old instructions are
//                retired from head.
//                
//                
//                
//  Create Date : original_time
//  Version     : v0.1 
//
//////////////////////////////////////////////////////////////////////////////////////////

module rob (


);




endmodule
